module test;


initial begin
    
end


jtkcpu_regs uut_regs (
    
);


endmodule